```vhdl
ENTITY error_example_solution IS
    PORT (
        clk : IN STD_LOGIC;
        rst : IN STD_LOGIC;
        data_in : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
        data_out : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END ENTITY error_example_solution;

ARCHITECTURE behavioral OF error_example_solution IS
    SIGNAL internal_data : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
BEGIN
    PROCESS (clk, rst, data_in) -- Corrected sensitivity list
    BEGIN
        IF rst = '1' THEN
            internal_data <= "00000000";
        ELSIF rising_edge(clk) THEN
            internal_data <= data_in;
        END IF;
    END PROCESS;

    data_out <= internal_data; 

END ARCHITECTURE behavioral;
```